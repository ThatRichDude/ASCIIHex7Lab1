/* Date: */
module sup(input A);
/* 
** Error: (vlog-13069) C:/Users/richardrojas/Dropbox (ASU)/Courses/Fall 2023/EEE 333/Lab/Lab One/ASCII_Code_All_RR.v(149): near "endmodule": syntax error, unexpected endmodule.

*/
endmodule;
